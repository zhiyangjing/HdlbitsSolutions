module top_module(output one);
    initial begin
        $display("asdf");
        $display("ssdf");
    end
endmodule


 
