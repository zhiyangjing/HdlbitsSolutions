module top_module( 
    input a, b, sel,
    output out ); 
  assign out = a & ~sel || b & sel;
endmodule
